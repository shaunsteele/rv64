// s_axi_lite_pkg.sv

`include "uvm_macros.svh"

package s_axi_lite_pkg;

import uvm_pkg::*;

`include "axi_lite_seq_item.sv"
`include "axi_lite_cfg.sv"
`include "s_axi_lite_monitor.sv"
`include "s_axi_lite_agent.sv"

endpackage
