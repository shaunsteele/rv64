// fetch_pkg.sv

`include "uvm_macros.svh"

package fetch_pkg;

import uvm_pkg::*;

`include "fetch_env.sv"
`include "fetch_base_test.sv"

endpackage
