// tb_store_pkg.sv

`include "uvm_macros.svh"

package tb_store_pkg;

import uvm_pkg::*;

`include "store_base_test.sv"

endpackage
